library verilog;
use verilog.vl_types.all;
entity Carry_Lookahead_32bits_vlg_vec_tst is
end Carry_Lookahead_32bits_vlg_vec_tst;
