library verilog;
use verilog.vl_types.all;
entity ripple_32_vlg_vec_tst is
end ripple_32_vlg_vec_tst;
